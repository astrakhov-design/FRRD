package tb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "tb_test.sv"

endpackage